module top(
	);
	
endmodule