//main decode
`define R_TYPE 	6'b000000
`define LW 		6'b100011
`define SW 		6'b101011
`define BEQ 	6'b000100
`define ADDI 	6'b001000
`define J 		6'b000010